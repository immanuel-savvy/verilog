module simple_function ();

function my_function;
input a,b,c,d;
  begin
    my_function = ((a+b) + (c-d));
  end
endfunction

endmodule // simple_function