module arithmetic_operators();

initial begin
  $display("5 + 10 = %d", 5 + 10);
  $display("5 - 10 = %d", 5 - 10);
  $display("10 - 5 = %d", 10 - 5);
  $display("5 * 10 = %d", 5 * 10);
  $display("10 / 5 = %d", 10 / 5);
  $display("10 %s 3 = %d",);
  $display("+5 = %d", +5);
  $display("-5 = %d", -5);
  #10 $finish;
end

endmodule